`timescale 1 ns / 10 ps
module cos_tb();
  // ----------------------------------
  // 參數與訊號宣告
  // ----------------------------------
  localparam T = 20;             // 時脈週期 (20 ns)
  reg clk;                       // 時脈訊號
  reg [5:0] addr;                // 輸入位址（假設最多64個資料點）
  wire [4:0] data;               // 從 sin 模組輸出的資料

  // ----------------------------------
  // DUT 實例化（Design Under Test）
  // ----------------------------------
  cos uut (
    .clk(clk),
    .addr(addr),
    .data(data)
  );

  // ----------------------------------
  // 時脈產生器：20ns 週期，50% duty cycle
  // ----------------------------------
  always begin
    clk = 1'b1;
    #(T / 2);
    clk = 1'b0;
    #(T / 2);
  end

  // ----------------------------------
  // 位址遞增：每個負緣時，addr + 1
  // ----------------------------------
  always @(negedge clk) begin
    addr <= addr + 1'b1;
  end

  // ----------------------------------
  // 初始條件與模擬結束控制
  // ----------------------------------
  initial begin
    addr = 6'b000000;         // 初始位址為 0
    #(128 * T);               // 模擬 128 個時脈週期
    $stop;                    // 結束模擬
  end

endmodule
